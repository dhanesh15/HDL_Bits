//Link : https://hdlbits.01xz.net/wiki/Zero
//Explanation: Output must be constant 0

module top_module(
    output zero
);// Module body starts after semicolon
	assign zero = 0;
endmodule
