//Link : https://hdlbits.01xz.net/wiki/Step_one
//Explanation: The expectation is to drive 1 to the output

module top_module( output one );

// Insert your code here
    assign one = 1;

endmodule
