//Link : https://hdlbits.01xz.net/wiki/Wire
//Explanation : Expected module should work like a wire

module top_module( input in, output out );
	assign out = in;
endmodule
