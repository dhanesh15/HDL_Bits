//Link : https://hdlbits.01xz.net/wiki/Exams/m2014_q4h
//Explanation : Output should be equal to the input

module top_module (
    input in,
    output out);
    
    assign out = in;

endmodule
