//Link : https://hdlbits.01xz.net/wiki/Sim/circuit1
//Explanation : Output is 1 when both inputs are 1, this resembles AND Gate

module top_module (
    input a,
    input b,
    output q );//

    assign q = a & b; // Fix me

endmodule
