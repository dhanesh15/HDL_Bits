//Link : https://hdlbits.01xz.net/wiki/Exams/m2014_q4i
//Explanation : Output should be tied to GND (or 0)

module top_module (
    output out);
    assign out = 1'b0;
endmodule
