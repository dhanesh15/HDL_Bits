//Link: https://hdlbits.01xz.net/wiki/Notgate
//Explanation: Module should work like a NOT Gate

module top_module( input in, output out );
    not (out , in );
endmodule
