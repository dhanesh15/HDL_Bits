//Link : https://hdlbits.01xz.net/wiki/Andgate
//Explanation : Module should work like an AND Gate

module top_module( 
    input a, 
    input b, 
    output out );
    assign out = a & b;

endmodule
